class i2c_master_transaction;
//TODO:
endclass